`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.02.2018 13:06:06
// Design Name: 
// Module Name: read_input_bram
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*
module read_input_bram(
input clk,
input reset,
input en,
input [17:0] addr,
output [15:0] data
    );

reg  
 input BRAM_PORTA_clk;
 input [15:0]BRAM_PORTA_din;
 input BRAM_PORTA_en;
 input [1:0]BRAM_PORTA_we;
 input [17:0]BRAM_PORTB_addr;
 input BRAM_PORTB_clk;
 output [15:0]BRAM_PORTB_dout;
 input BRAM_PORTB_en;
 input_bram bram
       (.BRAM_PORTA_addr(addr),
        .BRAM_PORTA_clk(clk),
        .BRAM_PORTA_en(en),
        .BRAM_PORTA_we(,
        .BRAM_PORTB_addr,
        .BRAM_PORTB_clk,
        .BRAM_PORTB_dout,
        .BRAM_PORTB_en);
    
endmodule
*/